//-----------------------------------------------------------------------------
//
// Title       : dispense
// Design      : DSD_Project
// Author      : shimu
// Company     : hp
//
//-----------------------------------------------------------------------------
//
// File        : C:/Users/HP/Downloads/DSD_Project/DSD_Project/DSD_Project/src/dispense.v
// Generated   : Mon Jan 20 01:30:38 2025
// From        : Interface description file
// By          : ItfToHdl ver. 1.0
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps

//{{ Section below this comment is automatically maintained
//    and may be overwritten
//{module {dispense}}

module dispense ( C ,En ,O );

input C;
wire C;
input En;
wire En;
output O;
wire O;


assign O = C & En;

//}} End of automatically maintained section

// Enter your statements here //

endmodule
